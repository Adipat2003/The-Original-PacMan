module map_font_rom(
    input [4:0] addr,
    output [15:0] data				 
);

	parameter ADDR_WIDTH = 5;
	parameter DATA_WIDTH = 16;
	
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = {
	    // Fill   
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        16'b0000000000000000,
        // No Fill
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111,
        16'b1111111111111111
	};
    
    assign data = ROM[addr];
    
endmodule
