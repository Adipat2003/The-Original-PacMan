module scared_ghost (
	input logic [7:0] address,
	output logic [3:0] q
);

logic [3:0] memory [0:255] /* synthesis ram_init_file = "./pac/pac.COE" */;

always_comb 
begin
	q = memory[address];
end

always_comb
begin
    memory [0] = 4'h1;
    memory [1] = 4'h1;
    memory [2] = 4'h1;
    memory [3] = 4'h1;
    memory [4] = 4'h1;
    memory [5] = 4'h1;
    memory [6] = 4'h1;
    memory [7] = 4'h1;
    memory [8] = 4'h1;
    memory [9] = 4'h1;
    memory [10] = 4'h1;
    memory [11] = 4'h1;
    memory [12] = 4'h1;
    memory [13] = 4'h1;
    memory [14] = 4'h1;
    memory [15] = 4'h1;
    memory [16] = 4'h1;
    memory [17] = 4'h1;
    memory [18] = 4'h1;
    memory [19] = 4'h1;
    memory [20] = 4'h1;
    memory [21] = 4'h1;
    memory [22] = 4'h0;
    memory [23] = 4'h0;
    memory [24] = 4'h0;
    memory [25] = 4'h0;
    memory [26] = 4'h1;
    memory [27] = 4'h1;
    memory [28] = 4'h1;
    memory [29] = 4'h1;
    memory [30] = 4'h1;
    memory [31] = 4'h1;
    memory [32] = 4'h1;
    memory [33] = 4'h1;
    memory [34] = 4'h1;
    memory [35] = 4'h1;
    memory [36] = 4'h0;
    memory [37] = 4'h0;
    memory [38] = 4'h0;
    memory [39] = 4'h0;
    memory [40] = 4'h0;
    memory [41] = 4'h0;
    memory [42] = 4'h0;
    memory [43] = 4'h0;
    memory [44] = 4'h1;
    memory [45] = 4'h1;
    memory [46] = 4'h1;
    memory [47] = 4'h1;
    memory [48] = 4'h1;
    memory [49] = 4'h1;
    memory [50] = 4'h1;
    memory [51] = 4'h0;
    memory [52] = 4'h0;
    memory [53] = 4'h0;
    memory [54] = 4'h0;
    memory [55] = 4'h0;
    memory [56] = 4'h0;
    memory [57] = 4'h0;
    memory [58] = 4'h0;
    memory [59] = 4'h0;
    memory [60] = 4'h0;
    memory [61] = 4'h1;
    memory [62] = 4'h1;
    memory [63] = 4'h1;
    memory [64] = 4'h1;
    memory [65] = 4'h1;
    memory [66] = 4'h0;
    memory [67] = 4'h0;
    memory [68] = 4'h0;
    memory [69] = 4'h0;
    memory [70] = 4'h0;
    memory [71] = 4'h0;
    memory [72] = 4'h0;
    memory [73] = 4'h0;
    memory [74] = 4'h0;
    memory [75] = 4'h0;
    memory [76] = 4'h0;
    memory [77] = 4'h0;
    memory [78] = 4'h1;
    memory [79] = 4'h1;
    memory [80] = 4'h1;
    memory [81] = 4'h1;
    memory [82] = 4'h0;
    memory [83] = 4'h0;
    memory [84] = 4'h0;
    memory [85] = 4'h0;
    memory [86] = 4'h0;
    memory [87] = 4'h0;
    memory [88] = 4'h0;
    memory [89] = 4'h0;
    memory [90] = 4'h0;
    memory [91] = 4'h0;
    memory [92] = 4'h0;
    memory [93] = 4'h0;
    memory [94] = 4'h1;
    memory [95] = 4'h1;
    memory [96] = 4'h1;
    memory [97] = 4'h1;
    memory [98] = 4'h0;
    memory [99] = 4'h0;
    memory [100] = 4'h0;
    memory [101] = 4'h2;
    memory [102] = 4'h2;
    memory [103] = 4'h0;
    memory [104] = 4'h0;
    memory [105] = 4'h2;
    memory [106] = 4'h2;
    memory [107] = 4'h0;
    memory [108] = 4'h0;
    memory [109] = 4'h0;
    memory [110] = 4'h1;
    memory [111] = 4'h1;
    memory [112] = 4'h1;
    memory [113] = 4'h0;
    memory [114] = 4'h0;
    memory [115] = 4'h0;
    memory [116] = 4'h0;
    memory [117] = 4'h2;
    memory [118] = 4'h2;
    memory [119] = 4'h0;
    memory [120] = 4'h0;
    memory [121] = 4'h2;
    memory [122] = 4'h2;
    memory [123] = 4'h0;
    memory [124] = 4'h0;
    memory [125] = 4'h0;
    memory [126] = 4'h0;
    memory [127] = 4'h1;
    memory [128] = 4'h1;
    memory [129] = 4'h0;
    memory [130] = 4'h0;
    memory [131] = 4'h0;
    memory [132] = 4'h0;
    memory [133] = 4'h0;
    memory [134] = 4'h0;
    memory [135] = 4'h0;
    memory [136] = 4'h0;
    memory [137] = 4'h0;
    memory [138] = 4'h0;
    memory [139] = 4'h0;
    memory [140] = 4'h0;
    memory [141] = 4'h0;
    memory [142] = 4'h0;
    memory [143] = 4'h1;
    memory [144] = 4'h1;
    memory [145] = 4'h0;
    memory [146] = 4'h0;
    memory [147] = 4'h0;
    memory [148] = 4'h0;
    memory [149] = 4'h0;
    memory [150] = 4'h0;
    memory [151] = 4'h0;
    memory [152] = 4'h0;
    memory [153] = 4'h0;
    memory [154] = 4'h0;
    memory [155] = 4'h0;
    memory [156] = 4'h0;
    memory [157] = 4'h0;
    memory [158] = 4'h0;
    memory [159] = 4'h1;
    memory [160] = 4'h1;
    memory [161] = 4'h0;
    memory [162] = 4'h0;
    memory [163] = 4'h2;
    memory [164] = 4'h2;
    memory [165] = 4'h0;
    memory [166] = 4'h0;
    memory [167] = 4'h2;
    memory [168] = 4'h2;
    memory [169] = 4'h0;
    memory [170] = 4'h0;
    memory [171] = 4'h2;
    memory [172] = 4'h2;
    memory [173] = 4'h0;
    memory [174] = 4'h0;
    memory [175] = 4'h1;
    memory [176] = 4'h1;
    memory [177] = 4'h0;
    memory [178] = 4'h2;
    memory [179] = 4'h0;
    memory [180] = 4'h0;
    memory [181] = 4'h2;
    memory [182] = 4'h2;
    memory [183] = 4'h0;
    memory [184] = 4'h0;
    memory [185] = 4'h2;
    memory [186] = 4'h2;
    memory [187] = 4'h0;
    memory [188] = 4'h0;
    memory [189] = 4'h2;
    memory [190] = 4'h0;
    memory [191] = 4'h1;
    memory [192] = 4'h1;
    memory [193] = 4'h0;
    memory [194] = 4'h0;
    memory [195] = 4'h0;
    memory [196] = 4'h0;
    memory [197] = 4'h0;
    memory [198] = 4'h0;
    memory [199] = 4'h0;
    memory [200] = 4'h0;
    memory [201] = 4'h0;
    memory [202] = 4'h0;
    memory [203] = 4'h0;
    memory [204] = 4'h0;
    memory [205] = 4'h0;
    memory [206] = 4'h0;
    memory [207] = 4'h1;
    memory [208] = 4'h1;
    memory [209] = 4'h0;
    memory [210] = 4'h0;
    memory [211] = 4'h0;
    memory [212] = 4'h0;
    memory [213] = 4'h1;
    memory [214] = 4'h0;
    memory [215] = 4'h0;
    memory [216] = 4'h0;
    memory [217] = 4'h0;
    memory [218] = 4'h1;
    memory [219] = 4'h0;
    memory [220] = 4'h0;
    memory [221] = 4'h0;
    memory [222] = 4'h0;
    memory [223] = 4'h1;
    memory [224] = 4'h1;
    memory [225] = 4'h1;
    memory [226] = 4'h0;
    memory [227] = 4'h0;
    memory [228] = 4'h1;
    memory [229] = 4'h1;
    memory [230] = 4'h1;
    memory [231] = 4'h0;
    memory [232] = 4'h0;
    memory [233] = 4'h1;
    memory [234] = 4'h1;
    memory [235] = 4'h1;
    memory [236] = 4'h0;
    memory [237] = 4'h0;
    memory [238] = 4'h1;
    memory [239] = 4'h1;
    memory [240] = 4'h1;
    memory [241] = 4'h1;
    memory [242] = 4'h1;
    memory [243] = 4'h1;
    memory [244] = 4'h1;
    memory [245] = 4'h1;
    memory [246] = 4'h1;
    memory [247] = 4'h1;
    memory [248] = 4'h1;
    memory [249] = 4'h1;
    memory [250] = 4'h1;
    memory [251] = 4'h1;
    memory [252] = 4'h1;
    memory [253] = 4'h1;
    memory [254] = 4'h1;
    memory [255] = 4'h1;

end

endmodule
